0000011300000093
0000021300000193
0000031300000293
0000041300000393
0000051300000493
0000061300000593
0000071300000693
0000081300000793
0000091300000893
00000A1300000993
00000B1300000A93
00000C1300000B93
00000D1300000C93
00000E1300000D93
00000F1300000E93
FF09011700000F93
000011B7F8410113
0001A023403101B3
FE219CE300418193
0281819300000197
000A07B730519073
0FF0000F7C079073
0000006F068000EF
0000001300000013
00B12623FF010113
342025F300C12423
008126030005DA63
0101011300C12583
0081260330200073
0101011300C12583
00000000FC5FF06F
0000194100000000
0100766373697200
337672050000000F
0000003070326932
F8300713900007B7
0007842300E78C23
00E7802300E00713
0000001300000013
0030071300000013
0007842300E78C23
00E78823FC000713
0287478390000737
FE078CE30207F793
0210071328C00793
00E68023900006B7
001787930017C703
2C400593FE071AE3
900007372C900613
0287478300058693
FE078CE30017F793
0016869300074783
FEF68FA300178793
02874783FED612E3
FE078CE30207F793
FC0786E32C404783
00F7002300058693
001686930016C783
FB5FF06FFE079AE3
00112623FF010113
900007B7F39FF0EF
00E78C23F8300713
00E0071300078423
0000001300E78023
0000001300000013
00E78C2300300713
FC00071300078423
0000806700E78823
00078C6300054783
00F7002390000737
0015051300154783
00008067FE079AE3
0287478390000737
FE078CE30017F793
0FF5751300074503
9000073700008067
0207F79302874783
00054783FE078CE3
9000073700078C63
0015478300F70023
FE079AE300150513
7365742100008067
3A434347000A2A74
392029554E472820
001B4100302E322E
0076637369720000
0510040000001101
3070326932337672
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
