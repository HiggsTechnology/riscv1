0000011300000093
0000021300000193
0000031300000293
0000041300000393
0000051300000493
0000061300000593
0000071300000693
0000081300000793
0000091300000893
00000A1300000993
00000B1300000A93
00000C1300000B93
00000D1300000C93
00000E1300000D93
00000F1300000E93
FF09011700000F93
000011B7F8410113
0001A023403101B3
FE219CE300418193
0281819300000197
4080079330519073
000A07B77F97A073
0FF0000F7C079073
0000006F058000EF
00B12623FF010113
342025F300C12423
008126030005DA63
0101011300C12583
0081260330200073
0101011300C12583
00001941FCDFF06F
0100766373697200
337672050000000F
0000003070326932
0680071317000793
00E6A423900406B7
001787930017C703
19800793FE071AE3
900406B707400713
0017C70300E6A423
FE071AE300178793
000080670006A623
00078C6300054783
00F7242390040737
0015051300154783
00008067FE079AE3
6F77206F6C6C6568
696874202C646C72
6E75662073692073
6574206E6F697463
000000000A217473
6C69772074736574
697320646E65206C
6E6F6974616C756D
3A43434700000000
392029554E472820
001B4100302E322E
0076637369720000
0510040000001101
3070326932337672
0000000000000000
